module ADDER();

endmodule
