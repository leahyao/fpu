module ADDER();


endmodule
